/*

Copyright (c) 2016-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * Generic IDDR module
 */
module iddr #
(
    // target ("SIM", "GENERIC", "XILINX", "ALTERA")
    parameter TARGET = "GENERIC",
    // IODDR style ("IODDR", "IODDR2")
    // Use IODDR for Virtex-4, Virtex-5, Virtex-6, 7 Series, Ultrascale
    // Use IODDR2 for Spartan-6
    parameter IODDR_STYLE = "IODDR2",
    // Width of register in bits
    parameter WIDTH = 1,
    parameter INSERT_BUFFERS = "FALSE"
)
(
    input  wire             clk,
    input  wire             rst,
    input  wire             en, 
    input  wire             en_vtc,
    input  wire             inc,
    input  wire             load,
    input  wire [8:0]      cnt_value_in,
    output wire [(WIDTH*9)-1:0]      cnt_value_out,
    input  wire refclk,
    output wire             rdy_idelay,
    // Data input   

    input  wire [WIDTH-1:0] d,

    output wire [WIDTH-1:0] q1,
    output wire [WIDTH-1:0] q2
);

/*

Provides a consistent input DDR flip flop across multiple FPGA families
              _____       _____       _____       _____       ____
    clk  ____/     \_____/     \_____/     \_____/     \_____/
         _ _____ _____ _____ _____ _____ _____ _____ _____ _____ _
    d    _X_D0__X_D1__X_D2__X_D3__X_D4__X_D5__X_D6__X_D7__X_D8__X_
         _______ ___________ ___________ ___________ ___________ _
    q1   _______X___________X____D0_____X____D2_____X____D4_____X_
         _______ ___________ ___________ ___________ ___________ _
    q2   _______X___________X____D1_____X____D3_____X____D5_____X_

*/
wire [WIDTH-1:0] d_int;
wire [WIDTH-1:0] delayed_data_int;
reg en_ff,en_ff1;
always @(posedge clk) begin
    en_ff <= en;
    en_ff1 <= en_ff;    
end
genvar n;

generate

if (INSERT_BUFFERS == "TRUE") begin
    for (genvar i = 0; i < WIDTH; i=i+1) begin
        IBUF IBUF_inst (
        .I(d[i]),
        .O(d_int[i])
        );
    end
end else begin
    assign d_int = d;
end

IDELAYCTRL #(
    .SIM_DEVICE("ULTRASCALE")  // Set the device version for simulation functionality (ULTRASCALE)
)
IDELAYCTRL_rx_inst (
    .RDY(rdy_idelay),       // 1-bit output: Ready output
    .REFCLK(refclk), // 1-bit input: Reference clock input
    .RST(0)        // 1-bit input: Active-High reset input. Asynchronous assert, synchronous deassert to
                       // REFCLK.
);

for (n = 0; n < WIDTH; n = n + 1) begin : iddr
      
   IDELAYE3 #(
      .CASCADE("NONE"),          // Cascade setting (MASTER, NONE, SLAVE_END, SLAVE_MIDDLE)
      .DELAY_FORMAT("COUNT"),     // Units of the DELAY_VALUE (COUNT, TIME)
      .DELAY_SRC("IDATAIN"),     // Delay input (DATAIN, IDATAIN)
      .DELAY_TYPE("VARIABLE"),      // Set the type of tap delay line (FIXED, VARIABLE, VAR_LOAD)
      .DELAY_VALUE(9'h19),           // Input delay value setting
      .IS_CLK_INVERTED(1'b0),    // Optional inversion for CLK
      .IS_RST_INVERTED(1'b0),    // Optional inversion for RST
      .REFCLK_FREQUENCY(300.0),  // IDELAYCTRL clock input frequency in MHz (200.0-800.0)
      .SIM_DEVICE("ULTRASCALE_PLUS"), // Set the device version for simulation functionality (ULTRASCALE)
      .UPDATE_MODE("ASYNC")      // Determines when updates to the delay will take effect (ASYNC, MANUAL, SYNC)
   )
   IDELAYE3_inst (
      .CASC_OUT(),       // 1-bit output: Cascade delay output to ODELAY input cascade
      .CNTVALUEOUT(cnt_value_out[(n*9)+8 : n*9 ]), // 9-bit output: Counter value output
      .DATAOUT(delayed_data_int[n]),         // 1-bit output: Delayed data output
      .CASC_IN(0),         // 1-bit input: Cascade delay input from slave ODELAY CASCADE_OUT
      .CASC_RETURN(0), // 1-bit input: Cascade delay returning from slave ODELAY DATAOUT
      .CE(en_ff & ~en_ff1),                   // 1-bit input: Active-High enable increment/decrement input
      .CLK(clk),                 // 1-bit input: Clock input
      .CNTVALUEIN(cnt_value_in),   // 9-bit input: Counter value input
      .DATAIN(0),           // 1-bit input: Data input from the logic
      .EN_VTC(en_vtc),           // 1-bit input: Keep delay constant over VT
      .IDATAIN(d_int[n]),         // 1-bit input: Data input from the IOBUF
      .INC(inc),                 // 1-bit input: Increment / Decrement tap delay input
      .LOAD(load),               // 1-bit input: Load DELAY_VALUE input
      .RST(rst)                  // 1-bit input: Asynchronous Reset to the DELAY_VALUE
   );

end
    reg [WIDTH-1:0] d_reg_1 = {WIDTH{1'b0}};
    reg [WIDTH-1:0] d_reg_2 = {WIDTH{1'b0}};

    reg [WIDTH-1:0] q_reg_1 = {WIDTH{1'b0}};
    reg [WIDTH-1:0] q_reg_2 = {WIDTH{1'b0}};

    always @(negedge clk) begin
        d_reg_1 <= delayed_data_int;
    end

    always @(posedge clk) begin
        d_reg_2 <= delayed_data_int;
    end

    always @(posedge clk) begin
        q_reg_1 <= d_reg_1;
        q_reg_2 <= d_reg_2;
    end

    assign q1 = q_reg_1;
    assign q2 = q_reg_2;

endgenerate

endmodule

`resetall
