/*

Copyright (c) 2015-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * 1G Ethernet MAC with GMII interface
 */
module eth_mac_1g_gmii #
(
    // target ("SIM", "GENERIC", "XILINX", "ALTERA")
    parameter TARGET = "GENERIC",
    // IODDR style ("IODDR", "IODDR2")
    // Use IODDR for Virtex-4, Virtex-5, Virtex-6, 7 Series, Ultrascale
    // Use IODDR2 for Spartan-6
    parameter IODDR_STYLE = "IODDR2",
    // Clock input style ("BUFG", "BUFR", "BUFIO", "BUFIO2")
    // Use BUFR for Virtex-5, Virtex-6, 7-series
    // Use BUFG for Ultrascale
    // Use BUFIO2 for Spartan-6
    parameter CLOCK_INPUT_STYLE = "BUFIO2",
    parameter ENABLE_PADDING = 1,
    parameter MIN_FRAME_LENGTH = 64
)
(
    input  wire        gtx_clk,
    input  wire        gtx_rst,
    output wire        rx_clk,
    output wire        rx_rst,
    output wire        tx_clk,
    output wire        tx_rst,

    /*
     * AXI input
     */
    input  wire [7:0]  tx_axis_tdata,
    input  wire        tx_axis_tvalid,
    output wire        tx_axis_tready,
    input  wire        tx_axis_tlast,
    input  wire        tx_axis_tuser,

    /*
     * AXI output
     */
    output wire [7:0]  rx_axis_tdata,
    output wire        rx_axis_tvalid,
    output wire        rx_axis_tlast,
    output wire        rx_axis_tuser,

    /*
     * GMII interface
     */
    input  wire        gmii_rx_clk,
    input  wire [7:0]  gmii_rxd,
    input  wire        gmii_rx_dv,
    input  wire        gmii_rx_er,
    // debug output
    output  reg [7:0]  gmii_rxd_out,
    output  reg        gmii_rx_dv_out,
    output  reg        gmii_rx_er_out, 
    output reg [7:0]  mac_gmii_rxd_out,
    output reg       mac_gmii_rx_dv_out,
    output reg       mac_gmii_rx_er_out,


    output wire [2:0] state_reg_out,
    output wire [2:0] state_next_out,
    output wire reset_crc_out,
    output wire update_crc_out,
    
    output wire mii_odd_out,
    output wire in_frame_out,
    
    output wire [7:0] gmii_rxd_d0_out,
    output wire [7:0] gmii_rxd_d1_out,
    output wire [7:0] gmii_rxd_d2_out,
    output wire [7:0] gmii_rxd_d3_out,
    output wire [7:0] gmii_rxd_d4_out,
    
    output wire gmii_rx_dv_d0_out,
    output wire gmii_rx_dv_d1_out,
    output wire gmii_rx_dv_d2_out,
    output wire gmii_rx_dv_d3_out,
    output wire gmii_rx_dv_d4_out,
    
    output wire gmii_rx_er_d0_out,
    output wire gmii_rx_er_d1_out,
    output wire gmii_rx_er_d2_out,
    output wire gmii_rx_er_d3_out,
    output wire gmii_rx_er_d4_out,
    
    output wire [7:0] m_axis_tdata_reg_out,
    output wire [7:0] m_axis_tdata_next_out,
    output wire m_axis_tvalid_reg_out,
    output wire m_axis_tvalid_next_out,
    output wire m_axis_tlast_reg_out, 
    output wire m_axis_tlast_next_out,
    output wire m_axis_tuser_reg_out, 
    output wire m_axis_tuser_next_out,
    
    output wire start_packet_int_reg_out,
    output wire start_packet_reg_out,
    output wire error_bad_frame_reg_out, 
    output wire error_bad_frame_next_out,
    output wire error_bad_fcs_reg_out,
    output wire error_bad_fcs_next_out,
    
    output wire [31-1:0] ptp_ts_reg_out,
    
    output wire [31:0] crc_state_out,
    output wire [31:0] crc_next_out,

    output wire clk_enable_out,
    output wire mii_select_out,
    
    output wire cfg_rx_enable_out,   
   
    input  wire        mii_tx_clk,
    output wire        gmii_tx_clk,
    output wire [7:0]  gmii_txd,
    output wire        gmii_tx_en,
    output wire        gmii_tx_er,

    /*
     * Status
     */
    output wire        tx_error_underflow,
    output wire        rx_error_bad_frame,
    output wire        rx_error_bad_fcs,
    output wire [1:0]  speed,

    /*
     * Configuration
     */
    input  wire [7:0]  cfg_ifg,
    input  wire        cfg_tx_enable,
    input  wire        cfg_rx_enable
);

wire [7:0]  mac_gmii_rxd;
wire        mac_gmii_rx_dv;
wire        mac_gmii_rx_er;
wire [7:0]  mac_gmii_txd;
wire        mac_gmii_tx_en;
wire        mac_gmii_tx_er;
always @(posedge rx_clk) begin
    gmii_rxd_out<=gmii_rxd;
    gmii_rx_dv_out<=gmii_rx_dv;
    gmii_rx_er_out<=gmii_rx_er; 
    mac_gmii_rxd_out<=mac_gmii_rxd;
    mac_gmii_rx_dv_out<=mac_gmii_rx_dv;
    mac_gmii_rx_er_out<=mac_gmii_rx_er;
end

reg [1:0] speed_reg = 2'b10;
reg mii_select_reg = 1'b0;

(* srl_style = "register" *)
reg [1:0] tx_mii_select_sync = 2'd0;

always @(posedge tx_clk) begin
    tx_mii_select_sync <= {tx_mii_select_sync[0], mii_select_reg};
end

(* srl_style = "register" *)
reg [1:0] rx_mii_select_sync = 2'd0;

always @(posedge rx_clk) begin
    rx_mii_select_sync <= {rx_mii_select_sync[0], mii_select_reg};
end

// PHY speed detection
reg [2:0] rx_prescale = 3'd0;

always @(posedge rx_clk) begin
    rx_prescale <= rx_prescale + 3'd1;
end

(* srl_style = "register" *)
reg [2:0] rx_prescale_sync = 3'd0;

always @(posedge gtx_clk) begin
    rx_prescale_sync <= {rx_prescale_sync[1:0], rx_prescale[2]};
end

reg [6:0] rx_speed_count_1 = 0;
reg [1:0] rx_speed_count_2 = 0;

always @(posedge gtx_clk) begin
    if (gtx_rst) begin
        rx_speed_count_1 <= 0;
        rx_speed_count_2 <= 0;
        speed_reg <= 2'b10;
        mii_select_reg <= 1'b0;
    end else begin
        rx_speed_count_1 <= rx_speed_count_1 + 1;
        
        if (rx_prescale_sync[1] ^ rx_prescale_sync[2]) begin
            rx_speed_count_2 <= rx_speed_count_2 + 1;
        end

        if (&rx_speed_count_1) begin
            // reference count overflow - 10M
            rx_speed_count_1 <= 0;
            rx_speed_count_2 <= 0;
            speed_reg <= 2'b00;
            mii_select_reg <= 1'b1;
        end

        if (&rx_speed_count_2) begin
            // prescaled count overflow - 100M or 1000M
            rx_speed_count_1 <= 0;
            rx_speed_count_2 <= 0;
            if (rx_speed_count_1[6:5]) begin
                // large reference count - 100M
                speed_reg <= 2'b01;
                mii_select_reg <= 1'b1;
            end else begin
                // small reference count - 1000M
                speed_reg <= 2'b10;
                mii_select_reg <= 1'b0;
            end
        end
    end
end

assign speed = speed_reg;

gmii_phy_if #(
    .TARGET(TARGET),
    .IODDR_STYLE(IODDR_STYLE),
    .CLOCK_INPUT_STYLE(CLOCK_INPUT_STYLE)
)
gmii_phy_if_inst (
    .clk(gtx_clk),
    .rst(gtx_rst),

    .mac_gmii_rx_clk(rx_clk),
    .mac_gmii_rx_rst(rx_rst),
    .mac_gmii_rxd(mac_gmii_rxd),
    .mac_gmii_rx_dv(mac_gmii_rx_dv),
    .mac_gmii_rx_er(mac_gmii_rx_er),
    .mac_gmii_tx_clk(tx_clk),
    .mac_gmii_tx_rst(tx_rst),
    .mac_gmii_txd(mac_gmii_txd),
    .mac_gmii_tx_en(mac_gmii_tx_en),
    .mac_gmii_tx_er(mac_gmii_tx_er),

    .phy_gmii_rx_clk(gmii_rx_clk),
    .phy_gmii_rxd(gmii_rxd),
    .phy_gmii_rx_dv(gmii_rx_dv),
    .phy_gmii_rx_er(gmii_rx_er),
    .phy_mii_tx_clk(mii_tx_clk),
    .phy_gmii_tx_clk(gmii_tx_clk),
    .phy_gmii_txd(gmii_txd),
    .phy_gmii_tx_en(gmii_tx_en),
    .phy_gmii_tx_er(gmii_tx_er),

    .mii_select(mii_select_reg)

);

eth_mac_1g #(
    .ENABLE_PADDING(ENABLE_PADDING),
    .MIN_FRAME_LENGTH(MIN_FRAME_LENGTH)
)
eth_mac_1g_inst (
    .tx_clk(tx_clk),
    .tx_rst(tx_rst),
    .rx_clk(rx_clk),
    .rx_rst(rx_rst),
    .tx_axis_tdata(tx_axis_tdata),
    .tx_axis_tvalid(tx_axis_tvalid),
    .tx_axis_tready(tx_axis_tready),
    .tx_axis_tlast(tx_axis_tlast),
    .tx_axis_tuser(tx_axis_tuser),
    .rx_axis_tdata(rx_axis_tdata),
    .rx_axis_tvalid(rx_axis_tvalid),
    .rx_axis_tlast(rx_axis_tlast),
    .rx_axis_tuser(rx_axis_tuser),
    .gmii_rxd(mac_gmii_rxd),
    .gmii_rx_dv(mac_gmii_rx_dv),
    .gmii_rx_er(mac_gmii_rx_er),
    .gmii_txd(mac_gmii_txd),
    .gmii_tx_en(mac_gmii_tx_en),
    .gmii_tx_er(mac_gmii_tx_er),
    .rx_clk_enable(1'b1),
    .tx_clk_enable(1'b1),
    .rx_mii_select(rx_mii_select_sync[1]),
    .tx_mii_select(tx_mii_select_sync[1]),
    .tx_error_underflow(tx_error_underflow),
    .rx_error_bad_frame(rx_error_bad_frame),
    .rx_error_bad_fcs(rx_error_bad_fcs),
    .cfg_ifg(cfg_ifg),
    .cfg_tx_enable(cfg_tx_enable),
    .cfg_rx_enable(cfg_rx_enable),
    .state_reg_out(state_reg_out),
    .state_next_out(state_next_out),
    .reset_crc_out(reset_crc_out),
    .update_crc_out(update_crc_out),
    
    .mii_odd_out(mii_odd_out),
    .in_frame_out(in_frame_out),
    
    .gmii_rxd_d0_out(gmii_rxd_d0_out),
    .gmii_rxd_d1_out(gmii_rxd_d1_out),
    .gmii_rxd_d2_out(gmii_rxd_d2_out),
    .gmii_rxd_d3_out(gmii_rxd_d3_out),
    .gmii_rxd_d4_out(gmii_rxd_d4_out),
    
    .gmii_rx_dv_d0_out(gmii_rx_dv_d0_out),
    .gmii_rx_dv_d1_out(gmii_rx_dv_d1_out),
    .gmii_rx_dv_d2_out(gmii_rx_dv_d2_out),
    .gmii_rx_dv_d3_out(gmii_rx_dv_d3_out),
    .gmii_rx_dv_d4_out(gmii_rx_dv_d4_out),
    
    .gmii_rx_er_d0_out(gmii_rx_er_d0_out),
    .gmii_rx_er_d1_out(gmii_rx_er_d1_out),
    .gmii_rx_er_d2_out(gmii_rx_er_d2_out),
    .gmii_rx_er_d3_out(gmii_rx_er_d3_out),
    .gmii_rx_er_d4_out(gmii_rx_er_d4_out),
    
    .m_axis_tdata_reg_out(m_axis_tdata_reg_out),
    .m_axis_tdata_next_out(m_axis_tdata_next_out),
    .m_axis_tvalid_reg_out(m_axis_tvalid_reg_out),
    .m_axis_tvalid_next_out(m_axis_tvalid_next_out),
    .m_axis_tlast_reg_out(m_axis_tlast_reg_out), 
    .m_axis_tlast_next_out(m_axis_tlast_next_out),
    .m_axis_tuser_reg_out(m_axis_tuser_reg_out), 
    .m_axis_tuser_next_out(m_axis_tuser_next_out),
    
    .start_packet_int_reg_out(start_packet_int_reg_out),
    .start_packet_reg_out(start_packet_reg_out),
    .error_bad_frame_reg_out(error_bad_frame_reg_out), 
    .error_bad_frame_next_out(error_bad_frame_next_out),
    .error_bad_fcs_reg_out(error_bad_fcs_reg_out),
    .error_bad_fcs_next_out(error_bad_fcs_next_out),
    .ptp_ts_reg_out(ptp_ts_reg_out),
    .crc_state_out(crc_state_out),
    .crc_next_out(crc_next_out),
    .clk_enable_out(clk_enable_out),
    .mii_select_out(mii_select_out),
    .cfg_rx_enable_out(cfg_rx_enable_out)   
);

endmodule

`resetall
